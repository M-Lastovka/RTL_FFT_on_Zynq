`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/05/2023 03:18:15 PM
// Design Name: 
// Module Name: sim_pckg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: package defining functions and parameters for TB
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


package axi_stream_pckg;
import dnn_pckg::*;

//AXI SLAVE

parameter S_TDATA_WDT = 32; //generated by setup_dnn_proj.py, do not edit manually 
parameter S_TID_WDT = 2; //generated by setup_dnn_proj.py, do not edit manually 
parameter S_FIFO_SIZE = 16; //generated by setup_dnn_proj.py, do not edit manually 
parameter S_FIFO_ADDR_WDT = $clog2(S_FIFO_SIZE);
parameter S_IF_BUFFER_SIZE = VLW_WDT/S_TDATA_WDT;
parameter S_IF_ADDR_WDT = 16; //TODO: make this more robust

parameter WEIGHT_S_AXIS_ID = 1;
parameter BIAS_S_AXIS_ID = 2;
parameter INPUT_S_AXIS_ID = 3;

//AXI MASTER

parameter M_TDATA_WDT = 32; //generated by setup_dnn_proj.py, do not edit manually 
parameter M_TID_WDT = 2; //generated by setup_dnn_proj.py, do not edit manually 
parameter M_FIFO_SIZE = 16; //generated by setup_dnn_proj.py, do not edit manually 
parameter M_FIFO_ADDR_WDT = $clog2(S_FIFO_SIZE);
parameter M_IF_BUFFER_SIZE = VLW_WDT/M_TDATA_WDT;

parameter M_PACKET_CNT = OUTPUT_MEM_SIZE*(VLW_WDT/M_TDATA_WDT);
parameter M_FIFO_WR_FINAL = ((M_PACKET_CNT % M_FIFO_SIZE)-1) == -1 ? M_FIFO_SIZE-1 : ((M_PACKET_CNT % M_FIFO_SIZE)-1); //value at which the fifo_wr_ptr should stop

endpackage